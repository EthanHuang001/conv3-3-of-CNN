`timescale 1ns/1ps
module tb_conv3x3_simple;

    // ʱ�Ӻ͸�λ
    reg clk;
    reg rst_n;
    
    // ģ������
    reg data_in_valid;
    reg [7:0] data_in_0, data_in_1, data_in_2;
    reg [7:0] data_in_3, data_in_4, data_in_5;
    reg [7:0] data_in_6, data_in_7, data_in_8;
    reg weight_en;
    reg signed [7:0] bias_data;
    reg [71:0] weights_data;
    
    // ģ�����
    wire data_out_valid;
    wire signed [17:0] data_out;
    
    // ʵ��������ģ��
    conv3x3 dut (
        .clk(clk), .rst_n(rst_n),
        .data_in_valid(data_in_valid),
        .data_in_0(data_in_0), .data_in_1(data_in_1), .data_in_2(data_in_2),
        .data_in_3(data_in_3), .data_in_4(data_in_4), .data_in_5(data_in_5),
        .data_in_6(data_in_6), .data_in_7(data_in_7), .data_in_8(data_in_8),
        .weight_en(weight_en), .bias_data(bias_data), .weights_data(weights_data),
        .data_out_valid(data_out_valid), .data_out(data_out)
    );
    
    // ʱ������ (100MHz)
    always #5 clk = ~clk;
    
    // ������֡5x5����ͼ��
    reg [7:0] frame1 [0:24]; // 5x5 = 25�����أ���һά�����ʾ
    reg [7:0] frame2 [0:24];
    reg [7:0] frame3 [0:24];
    
    integer i, j;
    
    initial begin
        // ��ʼ�������ļ�
        $dumpfile("conv3x3.vcd");
        $dumpvars(0, tb_conv3x3_simple);
        
        // ��ʼ���ź�
        clk = 0; rst_n = 1; data_in_valid = 0;
        weight_en = 0; bias_data = 8'sh00; weights_data = 72'b0;
        
        // ���ɲ���ͼ��
        generate_test_images();
        
        // ��λ����
        #10 rst_n = 0; #20 rst_n = 1; #10;
        
        // ����Ȩ��
        load_weights();
        
        // ������֡ͼ��
        process_frame(1); // ֡1: ����ģʽ
        #100;
        process_frame(2); // ֡2: ����ģʽ
        #100;  
        process_frame(3); // ֡3: ����ͻ��
        #200;
        
        $display("�������");
        $finish;
    end
    
    // ���ɲ���ͼ������
    task generate_test_images;
    begin
        // ֡1: ��1��25�ĵ���ģʽ
        for (i = 0; i < 25; i = i + 1) begin
            frame1[i] = i + 1;
        end
        
        // ֡2: ����ģʽ (1��2����)
        for (i = 0; i < 5; i = i + 1) begin
            for (j = 0; j < 5; j = j + 1) begin
                frame2[i*5+j] = ((i + j) % 2) ? 8'd1 : 8'd2;
            end
        end
        
        // ֡3: ����Ϊ10����ԵΪ1
        for (i = 0; i < 5; i = i + 1) begin
            for (j = 0; j < 5; j = j + 1) begin
                if (i >= 1 && i <= 3 && j >= 1 && j <= 3) 
                    frame3[i*5+j] = 8'd10;
                else 
                    frame3[i*5+j] = 8'd1;
            end
        end
        
        $display("����ͼ���������");
    end
    endtask
    
    // ����Ȩ������
    task load_weights;
    begin
        @(posedge clk);
        weight_en = 1;
        // Ȩ��ģʽ: [[1,1,1], [1,2,1], [1,1,1]]
        weights_data = 72'h01_01_01_01_02_01_01_01_01;
        @(posedge clk);
        weight_en = 0;
        $display("Ȩ�ؼ������: %h", weights_data);
    end
    endtask
    
    // ����֡ͼ������ - �޸���İ汾
    task process_frame;
    input integer frame_num;
    integer row, col;
    reg [7:0] current_pixel;
    begin
        $display("��ʼ����֡ %0d", frame_num);
        
        // ����3x3���ڴ���5x5ͼ�� (����3x3=9�����)
        for (row = 0; row < 3; row = row + 1) begin
            for (col = 0; col < 3; col = col + 1) begin
                @(posedge clk);
                data_in_valid = 1;
                
                // ����֡��ѡ���Ӧ��ͼ������
                case(frame_num)
                    1: current_pixel = frame1[row*5+col];
                    2: current_pixel = frame2[row*5+col];
                    3: current_pixel = frame3[row*5+col];
                endcase
                
                // �ṩ��ǰ3x3��������
                data_in_0 = (frame_num == 1) ? frame1[(row+0)*5+(col+0)] : 
                            (frame_num == 2) ? frame2[(row+0)*5+(col+0)] : frame3[(row+0)*5+(col+0)];
                data_in_1 = (frame_num == 1) ? frame1[(row+0)*5+(col+1)] : 
                            (frame_num == 2) ? frame2[(row+0)*5+(col+1)] : frame3[(row+0)*5+(col+1)];
                data_in_2 = (frame_num == 1) ? frame1[(row+0)*5+(col+2)] : 
                            (frame_num == 2) ? frame2[(row+0)*5+(col+2)] : frame3[(row+0)*5+(col+2)];
                data_in_3 = (frame_num == 1) ? frame1[(row+1)*5+(col+0)] : 
                            (frame_num == 2) ? frame2[(row+1)*5+(col+0)] : frame3[(row+1)*5+(col+0)];
                data_in_4 = (frame_num == 1) ? frame1[(row+1)*5+(col+1)] : 
                            (frame_num == 2) ? frame2[(row+1)*5+(col+1)] : frame3[(row+1)*5+(col+1)];
                data_in_5 = (frame_num == 1) ? frame1[(row+1)*5+(col+2)] : 
                            (frame_num == 2) ? frame2[(row+1)*5+(col+2)] : frame3[(row+1)*5+(col+2)];
                data_in_6 = (frame_num == 1) ? frame1[(row+2)*5+(col+0)] : 
                            (frame_num == 2) ? frame2[(row+2)*5+(col+0)] : frame3[(row+2)*5+(col+0)];
                data_in_7 = (frame_num == 1) ? frame1[(row+2)*5+(col+1)] : 
                            (frame_num == 2) ? frame2[(row+2)*5+(col+1)] : frame3[(row+2)*5+(col+1)];
                data_in_8 = (frame_num == 1) ? frame1[(row+2)*5+(col+2)] : 
                            (frame_num == 2) ? frame2[(row+2)*5+(col+2)] : frame3[(row+2)*5+(col+2)];
                
                $display("ʱ��%t: ֡%0d ����(%0d,%0d) ��������=%0d", 
                         $time, frame_num, row, col, data_in_4);
            end
        end
        
        @(posedge clk);
        data_in_valid = 0; // ֡�������
        $display("֡ %0d �������", frame_num);
    end
    endtask
    
    // ������
    always @(posedge clk) begin
        if (data_out_valid) begin
            $display("ʱ��%t: ������ = %0d", $time, data_out);
        end
    end

endmodule