`timescale 1ns / 1ps

module conv3x3 (
    input               clk,                // ʱ���ź�
    input               rst_n,              // �첽��λ���͵�ƽ��Ч
    input               data_in_valid,      // ����������Ч�ź�
    input       [7:0]   data_in_0,          // 3x3������������ (�޷���)
    input       [7:0]   data_in_1,
    input       [7:0]   data_in_2,
    input       [7:0]   data_in_3,
    input       [7:0]   data_in_4,
    input       [7:0]   data_in_5,
    input       [7:0]   data_in_6,
    input       [7:0]   data_in_7,
    input       [7:0]   data_in_8,
    input               weight_en,          // Ȩ��ʹ���ź�
    input signed [7:0]  bias_data,          // ƫ�����ݣ��з��ţ�Q1.7��ʽ
    input       [71:0]  weights_data,      // 72λȨ�����ݣ��ֽ�Ϊ9��8λȨ��
    
    output reg          data_out_valid,     // ���������Ч�ź�
    output reg signed [17:0] data_out        // ��������18λ�з�����(Q1.17��ʽ)
);

// Ȩ�ؼĴ�������72λweights_data�ֽ����
reg signed [7:0] weight_00, weight_01, weight_02;
reg signed [7:0] weight_10, weight_11, weight_12;
reg signed [7:0] weight_20, weight_21, weight_22;

// ����������ˮ�߼Ĵ������޷���ת�з��ţ�
reg signed [8:0] data_in_0_signed, data_in_1_signed, data_in_2_signed;
reg signed [8:0] data_in_3_signed, data_in_4_signed, data_in_5_signed;
reg signed [8:0] data_in_6_signed, data_in_7_signed, data_in_8_signed;

// ��һ����ˮ�ߣ��˷����
reg signed [16:0] prod_00, prod_01, prod_02;
reg signed [16:0] prod_10, prod_11, prod_12;
reg signed [16:0] prod_20, prod_21, prod_22;

// �ڶ�����ˮ�ߣ�����ͽ��
reg signed [17:0] sum_row0, sum_row1, sum_row2;

// ��������ˮ�ߣ��ܺͼ��㣨����һ����ˮ�ߣ�
reg signed [17:0] sum_total;

// ��Ч�ź���ˮ�ߣ�����һ�������ļ���
reg valid_d1, valid_d2, valid_d3, valid_d4;  // ��� valid_d4


always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        weight_00 <= 8'sb0; weight_01 <= 8'sb0; weight_02 <= 8'sb0;
        weight_10 <= 8'sb0; weight_11 <= 8'sb0; weight_12 <= 8'sb0;
        weight_20 <= 8'sb0; weight_21 <= 8'sb0; weight_22 <= 8'sb0;
    end else if (weight_en) begin
        // ��72λweights_data�зֽ�9��8λȨ��
        weight_00 <= $signed(weights_data[7:0]);
        weight_01 <= $signed(weights_data[15:8]);
        weight_02 <= $signed(weights_data[23:16]);
        weight_10 <= $signed(weights_data[31:24]);
        weight_11 <= $signed(weights_data[39:32]);
        weight_12 <= $signed(weights_data[47:40]);
        weight_20 <= $signed(weights_data[55:48]);
        weight_21 <= $signed(weights_data[63:56]);
        weight_22 <= $signed(weights_data[71:64]);
    end
end


always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        data_in_0_signed <= 9'sb0; data_in_1_signed <= 9'sb0; data_in_2_signed <= 9'sb0;
        data_in_3_signed <= 9'sb0; data_in_4_signed <= 9'sb0; data_in_5_signed <= 9'sb0;
        data_in_6_signed <= 9'sb0; data_in_7_signed <= 9'sb0; data_in_8_signed <= 9'sb0;
        valid_d1 <= 1'b0;
    end else begin
        data_in_0_signed <= {1'b0, data_in_0};
        data_in_1_signed <= {1'b0, data_in_1};
        data_in_2_signed <= {1'b0, data_in_2};
        data_in_3_signed <= {1'b0, data_in_3};
        data_in_4_signed <= {1'b0, data_in_4};
        data_in_5_signed <= {1'b0, data_in_5};
        data_in_6_signed <= {1'b0, data_in_6};
        data_in_7_signed <= {1'b0, data_in_7};
        data_in_8_signed <= {1'b0, data_in_8};
        valid_d1 <= data_in_valid;
    end
end


always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        prod_00 <= 17'sb0; prod_01 <= 17'sb0; prod_02 <= 17'sb0;
        prod_10 <= 17'sb0; prod_11 <= 17'sb0; prod_12 <= 17'sb0;
        prod_20 <= 17'sb0; prod_21 <= 17'sb0; prod_22 <= 17'sb0;
        valid_d2 <= 1'b0;
    end else begin
        prod_00 <= data_in_0_signed * weight_00;
        prod_01 <= data_in_1_signed * weight_01;
        prod_02 <= data_in_2_signed * weight_02;
        prod_10 <= data_in_3_signed * weight_10;
        prod_11 <= data_in_4_signed * weight_11;
        prod_12 <= data_in_5_signed * weight_12;
        prod_20 <= data_in_6_signed * weight_20;
        prod_21 <= data_in_7_signed * weight_21;
        prod_22 <= data_in_8_signed * weight_22;
        valid_d2 <= valid_d1;
    end
end


always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        sum_row0 <= 18'sb0;
        sum_row1 <= 18'sb0;
        sum_row2 <= 18'sb0;
        valid_d3 <= 1'b0;
    end else begin
        sum_row0 <= prod_00 + prod_01 + prod_02;
        sum_row1 <= prod_10 + prod_11 + prod_12;
        sum_row2 <= prod_20 + prod_21 + prod_22;
        valid_d3 <= valid_d2;
    end
end

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        sum_total <= 18'sb0;
        valid_d4 <= 1'b0;  // ��ʼ����������Ч�źżĴ���
    end else begin
        // �������н�����ܺ�
        sum_total <= sum_row0 + sum_row1 + sum_row2;
        // ��Ч�ź��ӳ�һ��
        valid_d4 <= valid_d3;
    end
end


always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        data_out <= 18'sb0;
        data_out_valid <= 1'b0;
    end else begin
        // ����ƫ�ã�ƫ��ΪQ1.7��ʽ����Ҫ����10λ���룩
        data_out <= sum_total + ({{10{bias_data[7]}}, bias_data, 1'b0});
        // ��Ч�ź�������ͬ�����
        data_out_valid <= valid_d4;
    end
end

endmodule